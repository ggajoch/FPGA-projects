
module unnamed (
	acq_data_in,
	acq_trigger_in,
	acq_clk);	

	input	[9:0]	acq_data_in;
	input	[0:0]	acq_trigger_in;
	input		acq_clk;
endmodule
