-- unnamed.vhd

-- Generated using ACDS version 14.0 200 at 2014.10.16.22:43:23

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unnamed is
	port (
		acq_data_in    : in std_logic_vector(9 downto 0) := (others => '0'); --     tap.acq_data_in
		acq_trigger_in : in std_logic_vector(0 downto 0) := (others => '0'); --        .acq_trigger_in
		acq_clk        : in std_logic                    := '0'              -- acq_clk.clk
	);
end entity unnamed;

architecture rtl of unnamed is
	component sld_signaltap is
		generic (
			sld_data_bits               : integer := 1;
			sld_sample_depth            : integer := 128;
			sld_ram_block_type          : string  := "AUTO";
			sld_storage_qualifier_mode  : string  := "OFF";
			sld_trigger_bits            : integer := 1;
			sld_trigger_level           : integer := 1;
			sld_trigger_in_enabled      : boolean := false;
			sld_enable_advanced_trigger : boolean := false;
			sld_trigger_level_pipeline  : integer := 1;
			sld_node_info               : integer := 1076736;
			sld_node_crc_bits           : integer := 32;
			sld_node_crc_hiword         : integer := 12345;
			sld_node_crc_loword         : integer := 19899
		);
		port (
			acq_data_in    : in std_logic_vector(9 downto 0) := (others => 'X'); -- acq_data_in
			acq_trigger_in : in std_logic_vector(0 downto 0) := (others => 'X'); -- acq_trigger_in
			acq_clk        : in std_logic                    := 'X'              -- clk
		);
	end component sld_signaltap;

begin

	signaltap_ii_logic_analyzer_0 : component sld_signaltap
		generic map (
			sld_data_bits               => 10,
			sld_sample_depth            => 128,
			sld_ram_block_type          => "AUTO",
			sld_storage_qualifier_mode  => "OFF",
			sld_trigger_bits            => 1,
			sld_trigger_level           => 1,
			sld_trigger_in_enabled      => false,
			sld_enable_advanced_trigger => false,
			sld_trigger_level_pipeline  => 1,
			sld_node_info               => 1076736,
			sld_node_crc_bits           => 32,
			sld_node_crc_hiword         => 39533,
			sld_node_crc_loword         => 62180
		)
		port map (
			acq_data_in    => acq_data_in,    --     tap.acq_data_in
			acq_trigger_in => acq_trigger_in, --        .acq_trigger_in
			acq_clk        => acq_clk         -- acq_clk.clk
		);

end architecture rtl; -- of unnamed
